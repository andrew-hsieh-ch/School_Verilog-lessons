module video (
    input clk,
    input reset_p,
    output reg [7:0]LED_ROW,
    output reg [7:0]LED1_ROW,
    output reg [7:0]LED2_ROW,
    output reg [7:0]LED_ROW3,
    output reg [7:0]LED_ROW4,
    output reg [7:0]LED_ROW5,
    output reg [7:0]LED_ROW6,
    output reg [7:0]LED_ROW7,
    output reg [7:0]LED_COL
);
    
localparam count_max = 25'd50000;

integer j;

reg [24:0] counter;

reg [7:0]map [167:0];
reg [7:0]map1[167:0];
reg [7:0]map2[167:0];
reg [7:0]map3[167:0];
reg [7:0]map4[167:0];
reg [7:0]map5[31:0];
reg [7:0]map6[31:0];
reg [7:0]map7[31:0];


reg [3:0]i;

wire time_flag;

assign time_flag = (counter == count_max - 1'b1) ? 1'b1 : 1'b0;

always @(posedge clk or posedge reset_p) begin
    if(reset_p)
        counter <= 25'd0;
    else
        counter <= (counter == count_max - 1'b1) ? 25'd0 : counter + 1'b1;
end

always @(posedge clk or posedge reset_p) begin
    if(reset_p)
        i <= 2'd0;
    else
        i <= (time_flag) ? i + 1'b1 : i;
end

always @(posedge clk or posedge reset_p) begin
    if(reset_p)
        LED_ROW <= 8'd0;
    else
        case (LED_COL)
            8'h01 : LED_ROW <= map[0 + {i,3'd0}] ; 
            8'h02 : LED_ROW <= map[1 + {i,3'd0}] ;
            8'h04 : LED_ROW <= map[2 + {i,3'd0}] ;
            8'h08 : LED_ROW <= map[3 + {i,3'd0}] ;
            8'h10 : LED_ROW <= map[4 + {i,3'd0}] ;
            8'h20 : LED_ROW <= map[5 + {i,3'd0}] ;
            8'h40 : LED_ROW <= map[6 + {i,3'd0}] ;
            8'h80 : LED_ROW <= map[7 + {i,3'd0}] ;
            default: LED_ROW <= 8'h00;
        endcase
end
always @(posedge clk or posedge reset_p) begin
    if(reset_p)
        LED1_ROW <= 8'd0;
    else
        case (LED_COL)
            8'h01 : LED1_ROW <= map1[0 + {i,3'd0}] ; 
            8'h02 : LED1_ROW <= map1[1 + {i,3'd0}] ;
            8'h04 : LED1_ROW <= map1[2 + {i,3'd0}] ;
            8'h08 : LED1_ROW <= map1[3 + {i,3'd0}] ;
            8'h10 : LED1_ROW <= map1[4 + {i,3'd0}] ;
            8'h20 : LED1_ROW <= map1[5 + {i,3'd0}] ;
            8'h40 : LED1_ROW <= map1[6 + {i,3'd0}] ;
            8'h80 : LED1_ROW <= map1[7 + {i,3'd0}] ;
            default: LED1_ROW <= 8'h00;
        endcase
end

always @(posedge clk or posedge reset_p) begin
    if(reset_p)
        LED2_ROW <= 8'd0;
    else
        case (LED_COL)
            8'h01 : LED2_ROW <= map2[0 + {i,3'd0}] ; 
            8'h02 : LED2_ROW <= map2[1 + {i,3'd0}] ;
            8'h04 : LED2_ROW <= map2[2 + {i,3'd0}] ;
            8'h08 : LED2_ROW <= map2[3 + {i,3'd0}] ;
            8'h10 : LED2_ROW <= map2[4 + {i,3'd0}] ;
            8'h20 : LED2_ROW <= map2[5 + {i,3'd0}] ;
            8'h40 : LED2_ROW <= map2[6 + {i,3'd0}] ;
            8'h80 : LED2_ROW <= map2[7 + {i,3'd0}] ;
            default: LED2_ROW <= 8'h00;
        endcase
end

always @(posedge clk or posedge reset_p) begin
    if(reset_p)
        LED_ROW3 <= 8'd0;
    else
        case (LED_COL)
            8'h01 : LED_ROW3 <= map3[0 + {i,3'd0}] ; 
            8'h02 : LED_ROW3 <= map3[1 + {i,3'd0}] ;
            8'h04 : LED_ROW3 <= map3[2 + {i,3'd0}] ;
            8'h08 : LED_ROW3 <= map3[3 + {i,3'd0}] ;
            8'h10 : LED_ROW3 <= map3[4 + {i,3'd0}] ;
            8'h20 : LED_ROW3 <= map3[5 + {i,3'd0}] ;
            8'h40 : LED_ROW3 <= map3[6 + {i,3'd0}] ;
            8'h80 : LED_ROW3 <= map3[7 + {i,3'd0}] ;
            default: LED_ROW3 <= 8'h00;
        endcase
end

always @(posedge clk or posedge reset_p) begin
    if(reset_p)
        LED_ROW4 <= 8'd0;
    else
        case (LED_COL)
            8'h01 : LED_ROW4 <= map4[0 + {i,3'd0}] ; 
            8'h02 : LED_ROW4 <= map4[1 + {i,3'd0}] ;
            8'h04 : LED_ROW4 <= map4[2 + {i,3'd0}] ;
            8'h08 : LED_ROW4 <= map4[3 + {i,3'd0}] ;
            8'h10 : LED_ROW4 <= map4[4 + {i,3'd0}] ;
            8'h20 : LED_ROW4 <= map4[5 + {i,3'd0}] ;
            8'h40 : LED_ROW4 <= map4[6 + {i,3'd0}] ;
            8'h80 : LED_ROW4 <= map4[7 + {i,3'd0}] ;
            default: LED_ROW4 <= 8'h00;
        endcase
end

always @(posedge clk or posedge reset_p) begin
    if(reset_p)
        LED_ROW5 <= 8'd0;
    else
        case (LED_COL)
            8'h01 : LED_ROW5 <= map5[0 + {i,3'd0}] ; 
            8'h02 : LED_ROW5 <= map5[1 + {i,3'd0}] ;
            8'h04 : LED_ROW5 <= map5[2 + {i,3'd0}] ;
            8'h08 : LED_ROW5 <= map5[3 + {i,3'd0}] ;
            8'h10 : LED_ROW5 <= map5[4 + {i,3'd0}] ;
            8'h20 : LED_ROW5 <= map5[5 + {i,3'd0}] ;
            8'h40 : LED_ROW5 <= map5[6 + {i,3'd0}] ;
            8'h80 : LED_ROW5 <= map5[7 + {i,3'd0}] ;
            default: LED_ROW5 <= 8'h00;
        endcase
end
always @(posedge clk or posedge reset_p) begin
    if(reset_p)
        LED_ROW6 <= 8'd0;
    else
        case (LED_COL)
            8'h01 : LED_ROW6 <= map6[0 + {i,3'd0}] ; 
            8'h02 : LED_ROW6 <= map6[1 + {i,3'd0}] ;
            8'h04 : LED_ROW6 <= map6[2 + {i,3'd0}] ;
            8'h08 : LED_ROW6 <= map6[3 + {i,3'd0}] ;
            8'h10 : LED_ROW6 <= map6[4 + {i,3'd0}] ;
            8'h20 : LED_ROW6 <= map6[5 + {i,3'd0}] ;
            8'h40 : LED_ROW6 <= map6[6 + {i,3'd0}] ;
            8'h80 : LED_ROW6 <= map6[7 + {i,3'd0}] ;
            default: LED_ROW6 <= 8'h00;
        endcase
end
always @(posedge clk or posedge reset_p) begin
    if(reset_p)
        LED_ROW7 <= 8'd0;
    else
        case (LED_COL)
            8'h01 : LED_ROW7 <= map7[0 + {i,3'd0}] ; 
            8'h02 : LED_ROW7 <= map7[1 + {i,3'd0}] ;
            8'h04 : LED_ROW7 <= map7[2 + {i,3'd0}] ;
            8'h08 : LED_ROW7 <= map7[3 + {i,3'd0}] ;
            8'h10 : LED_ROW7 <= map7[4 + {i,3'd0}] ;
            8'h20 : LED_ROW7 <= map7[5 + {i,3'd0}] ;
            8'h40 : LED_ROW7 <= map7[6 + {i,3'd0}] ;
            8'h80 : LED_ROW7 <= map7[7 + {i,3'd0}] ;
            default: LED_ROW7 <= 8'h00;
        endcase
end
always @(posedge clk or posedge reset_p) begin
    if(reset_p)
        LED_COL <= 8'h01;
    else
        LED_COL <= (LED_COL == 8'h80) ? 8'h01 : 
        {LED_COL[6:0],1'b0};
end

always @(posedge clk or posedge reset_p) begin
    if(reset_p)
    begin
        map[0] = 8'b00000000;//1
        map[1] = 8'b00000000;
        map[2] = 8'b00000000;
        map[3] = 8'b00001110;
        map[4] = 8'b00011011;
        map[5] = 8'b00010001;
        map[6] = 8'b00010001;
        map[7] = 8'b00010001;

        map[8] = 8'b00000000;//2
        map[9] = 8'b00000000;
        map[10] = 8'b00000000;
        map[11] = 8'b00001110;
        map[12] = 8'b00011011;
        map[13] = 8'b00010001;
        map[14] = 8'b00010001;
        map[15] = 8'b00010001;

        map[16] = 8'b00000000;//3
        map[17] = 8'b00000000;
        map[18] = 8'b00000000;
        map[19] = 8'b00001110;
        map[20] = 8'b00011011;
        map[21] = 8'b00010001;
        map[22] = 8'b00010001;
        map[23] = 8'b00010001;

        map[24] = 8'b00000000;//4
        map[25] = 8'b00000000;
        map[26] = 8'b00000000;
        map[27] = 8'b00001110;
        map[28] = 8'b00011011;
        map[29] = 8'b00010001;
        map[30] = 8'b00010001;
        map[31] = 8'b00010001;

		map[32] = 8'b00000000;//5
        map[33] = 8'b00000000;
        map[34] = 8'b00000000;
        map[35] = 8'b00001110;
        map[36] = 8'b00011011;
        map[37] = 8'b00010001;
        map[38] = 8'b00010001;
        map[39] = 8'b00010001;
        
        map[40] = 8'b00000000;//6
        map[41] = 8'b00000000;
        map[42] = 8'b00001110;
        map[43] = 8'b00001110;
        map[44] = 8'b00011011;
        map[45] = 8'b00010001;
        map[46] = 8'b00010001;
        map[47] = 8'b00010001;
        
        map[48] = 8'b00000000;//7
        map[49] = 8'b00000000;
        map[50] = 8'b00000000;
        map[51] = 8'b00001110;
        map[52] = 8'b00011011;
        map[53] = 8'b00010001;
        map[54] = 8'b00010001;
        map[55] = 8'b00010001;
        
        map[56] = 8'b00000000;//8
        map[57] = 8'b00000000;
        map[58] = 8'b00000000;
        map[59] = 8'b00001110;
        map[60] = 8'b00011011;
        map[61] = 8'b00010001;
        map[62] = 8'b00010001;
        map[63] = 8'b00010001;
        
        map[64] = 8'b00000000;//9
        map[65] = 8'b00000000;
        map[66] = 8'b00000000;
        map[67] = 8'b00001110;
        map[68] = 8'b00011011;
        map[69] = 8'b00010001;
        map[70] = 8'b00010001;
        map[71] = 8'b00010001;
        
        map[72] = 8'b00000000;//10
        map[73] = 8'b00000000;
        map[74] = 8'b00000000;
        map[75] = 8'b00001110;
        map[76] = 8'b00011011;
        map[77] = 8'b00010001;
        map[78] = 8'b00010001;
        map[79] = 8'b00010001;
        
        map[80] = 8'b00000000;//11
        map[81] = 8'b00000000;
        map[82] = 8'b00000000;
        map[83] = 8'b00001110;
        map[84] = 8'b00011011;
        map[85] = 8'b00010001;
        map[86] = 8'b00010001;
        map[87] = 8'b00010001;
        
        map[88] = 8'b00000000;//12
        map[89] = 8'b00000000;
        map[90] = 8'b00000000;
        map[91] = 8'b00001110;
        map[92] = 8'b00011011;
        map[93] = 8'b00010001;
        map[94] = 8'b00010001;
        map[95] = 8'b00010001;
       
        map[96] = 8'b00000000;//13
        map[97] = 8'b00000000;
        map[98] = 8'b00000000;
        map[99] = 8'b00001110;
        map[100] = 8'b00011011;
        map[101] = 8'b00100001;
        map[102] = 8'b00110001;
        map[103] = 8'b00010001;
        
        map[104] = 8'b00000000;//14
        map[105] = 8'b00000000;
        map[106] = 8'b00000000;
        map[107] = 8'b00001110;
        map[108] = 8'b00011011;
        map[109] = 8'b00100001;
        map[110] = 8'b00110001;
        map[111] = 8'b00010001;
        
        map[112] = 8'b00000000;//15
        map[113] = 8'b00000000;
        map[114] = 8'b00000000;
        map[115] = 8'b00001110;
        map[116] = 8'b00011011;
        map[117] = 8'b00100001;
        map[118] = 8'b00110001;
        map[119] = 8'b00010001;
        
        map[120] = 8'b00000000;//16
        map[121] = 8'b00000000;
        map[122] = 8'b00000000;
        map[123] = 8'b00001110;
        map[124] = 8'b00011011;
        map[125] = 8'b00100001;
        map[126] = 8'b00110001;
        map[127] = 8'b00010001;
        
        map[128] = 8'b00000000;//17
        map[129] = 8'b00000000;
        map[130] = 8'b00000000;
        map[131] = 8'b00001110;
        map[132] = 8'b00011011;
        map[133] = 8'b00100001;
        map[134] = 8'b00110001;
        map[135] = 8'b00010001;
        
        map[136] = 8'b00000000;//18
        map[137] = 8'b00000000;
        map[138] = 8'b00000111;
        map[139] = 8'b00001101;
        map[140] = 8'b00010000;
        map[141] = 8'b00011000;
        map[142] = 8'b00001000;
        map[143] = 8'b00001101;
        
        map[144] = 8'b00000000;//19
        map[145] = 8'b00000000;
        map[146] = 8'b00000011;
        map[147] = 8'b00000110;
        map[148] = 8'b00001000;
        map[149] = 8'b00001100;
        map[150] = 8'b00000100;
        map[151] = 8'b00000110;
        
        map[152] = 8'b00000000;//20
        map[153] = 8'b00000000;
        map[154] = 8'b00000000;
        map[155] = 8'b00000001;
        map[156] = 8'b00000010;
        map[157] = 8'b00000011;
        map[158] = 8'b00000001;
        map[159] = 8'b00000001;
        
        map[160] = 8'b00000000;//21
        map[161] = 8'b00000000;
        map[162] = 8'b00000000;
        map[163] = 8'b00000001;
        map[164] = 8'b00000010;
        map[165] = 8'b00000011;
        map[166] = 8'b00000001;
        map[167] = 8'b00000001;
        
    end
    else
        for(j = 0;j < 168;j = j + 1)
            map[j] = map[j];
end

always @(posedge clk or posedge reset_p) begin
    if(reset_p)
    begin
        map1[0] = 8'b00001010;//1
        map1[1] = 8'b00000100;
        map1[2] = 8'b00001110;
        map1[3] = 8'b00010101;
        map1[4] = 8'b00100100;
        map1[5] = 8'b00001010;
        map1[6] = 8'b00001010;
        map1[7] = 8'b00010001;

        map1[8] = 8'b00001010;//2
        map1[9] = 8'b00001110;
        map1[10] = 8'b00010101;
        map1[11] = 8'b00100100;
        map1[12] = 8'b00000100;
        map1[13] = 8'b00001010;
        map1[14] = 8'b00001010;
        map1[15] = 8'b00010001;

        map1[16] = 8'b00001010;//3
        map1[17] = 8'b00000100;
        map1[18] = 8'b00001110;
        map1[19] = 8'b00010101;
        map1[20] = 8'b00100100;
        map1[21] = 8'b00001010;
        map1[22] = 8'b00001010;
        map1[23] = 8'b00010001;

        map1[24] = 8'b00001010;//4
        map1[25] = 8'b00001110;
        map1[26] = 8'b00010101;
        map1[27] = 8'b00100100;
        map1[28] = 8'b00000100;
        map1[29] = 8'b00001010;
        map1[30] = 8'b00001010;
        map1[31] = 8'b00010001;
        
        map1[32] = 8'b00001010;//5
        map1[33] = 8'b00001110;
        map1[34] = 8'b00010101;
        map1[35] = 8'b00100100;
        map1[36] = 8'b00000100;
        map1[37] = 8'b00001010;
        map1[38] = 8'b00001010;
        map1[39] = 8'b00010001;
        
        map1[40] = 8'b00001010;//6
        map1[41] = 8'b00001110;
        map1[42] = 8'b00010101;
        map1[43] = 8'b00100100;
        map1[44] = 8'b00000100;
        map1[45] = 8'b00001010;
        map1[46] = 8'b00001010;
        map1[47] = 8'b00010001;
        
        map1[48] = 8'b00001010;//7
        map1[49] = 8'b00001110;
        map1[50] = 8'b00010101;
        map1[51] = 8'b00100100;
        map1[52] = 8'b00000100;
        map1[53] = 8'b00001010;
        map1[54] = 8'b00001010;
        map1[55] = 8'b00010001;
        
        map1[56] = 8'b00001010;//8
        map1[57] = 8'b00001110;
        map1[58] = 8'b00010101;
        map1[59] = 8'b00100100;
        map1[60] = 8'b00000100;
        map1[61] = 8'b00001010;
        map1[62] = 8'b00001010;
        map1[63] = 8'b00010001;
        
        map1[64] = 8'b00001010;//9
        map1[65] = 8'b00001110;
        map1[66] = 8'b00010101;
        map1[67] = 8'b00100100;
        map1[68] = 8'b00000100;
        map1[69] = 8'b00001010;
        map1[70] = 8'b00001010;
        map1[71] = 8'b00010001;
        
        map1[72] = 8'b00001010;//10
        map1[73] = 8'b00001110;
        map1[74] = 8'b00010101;
        map1[75] = 8'b00100100;
        map1[76] = 8'b00000100;
        map1[77] = 8'b00001010;
        map1[78] = 8'b00001010;
        map1[79] = 8'b00010001;
        
        map1[80] = 8'b00001010;//11
        map1[81] = 8'b00001110;
        map1[82] = 8'b00010101;
        map1[83] = 8'b00100100;
        map1[84] = 8'b00000100;
        map1[85] = 8'b00001010;
        map1[86] = 8'b00001010;
        map1[87] = 8'b00010001;
        
        map1[88] = 8'b00001010;//12
        map1[89] = 8'b00001110;
        map1[90] = 8'b00010101;
        map1[91] = 8'b00100100;
        map1[92] = 8'b00000100;
        map1[93] = 8'b00001010;
        map1[94] = 8'b00001010;
        map1[95] = 8'b00010001;
       
        map1[96] = 8'b00011010;//13
        map1[97] = 8'b00000100;
        map1[98] = 8'b00001111;
        map1[99] = 8'b00010100;
        map1[100] = 8'b00011110;
        map1[101] = 8'b000001001;
        map1[102] = 8'b00001000;
        map1[103] = 8'b00010000;
        
        map1[104] = 8'b00011010;//14
        map1[105] = 8'b00000101;
        map1[106] = 8'b00001110;
        map1[107] = 8'b00010100;
        map1[108] = 8'b00001110;
        map1[109] = 8'b00001001;
        map1[110] = 8'b00010000;
        map1[111] = 8'b00100000;
        
        map1[112] = 8'b00011010;//15
        map1[113] = 8'b00000101;
        map1[114] = 8'b00001110;
        map1[115] = 8'b00010100;
        map1[116] = 8'b00011110;
        map1[117] = 8'b00001001;
        map1[118] = 8'b00010000;
        map1[119] = 8'b00100000;
        
        map1[120] = 8'b00011010;//16
        map1[121] = 8'b00000100;
        map1[122] = 8'b00001111;
        map1[123] = 8'b00010100;
        map1[124] = 8'b00101110;
        map1[125] = 8'b00001001;
        map1[126] = 8'b00011000;
        map1[127] = 8'b00100000;
        
        map1[128] = 8'b00011010;//17
        map1[129] = 8'b00000100;
        map1[130] = 8'b00001111;
        map1[131] = 8'b00010100;
        map1[132] = 8'b00101110;
        map1[133] = 8'b00001001;
        map1[134] = 8'b00010000;
        map1[135] = 8'b00100000;
        
        map1[136] = 8'b00000010;//18
        map1[137] = 8'b00000111;
        map1[138] = 8'b00001010;
        map1[139] = 8'b00010110;
        map1[140] = 8'b00001001;
        map1[141] = 8'b00010000;
        map1[142] = 8'b00100000;
        map1[143] = 8'b00000001;
        
        map1[144] = 8'b00000001;//19
        map1[145] = 8'b00000011;
        map1[146] = 8'b00000101;
        map1[147] = 8'b00001011;
        map1[148] = 8'b00000100;
        map1[149] = 8'b00001000;
        map1[150] = 8'b00010000;
        map1[151] = 8'b00000001;
        
        map1[152] = 8'b00000000;//20
        map1[153] = 8'b00000000;
        map1[154] = 8'b00000001;
        map1[155] = 8'b00000010;
        map1[156] = 8'b00000001;
        map1[157] = 8'b00000010;
        map1[158] = 8'b00000100;
        map1[159] = 8'b00000000;
        
        map1[160] = 8'b00000000;//21
        map1[161] = 8'b00000000;
        map1[162] = 8'b00000001;
        map1[163] = 8'b00000010;
        map1[164] = 8'b00000001;
        map1[165] = 8'b00000010;
        map1[166] = 8'b00000101;
        map1[167] = 8'b00000000;
    end
    else
        for(j = 0;j < 168 ;j = j + 1)
            map1[j] = map1[j];
end

always @(posedge clk or posedge reset_p) begin
    if(reset_p)
    begin
        map2[0] = 8'b00000000;//1
        map2[1] = 8'b00000000;
        map2[2] = 8'b00000000;
        map2[3] = 8'b00000000;
        map2[4] = 8'b00000000;
        map2[5] = 8'b00000000;
        map2[6] = 8'b00000000;
        map2[7] = 8'b00000000;

        map2[8] = 8'b00000000;//2
        map2[9] = 8'b00000000;
        map2[10] = 8'b00000000;
        map2[11] = 8'b00000000;
        map2[12] = 8'b00000000;
        map2[13] = 8'b00000000;
        map2[14] = 8'b00000000;
        map2[15] = 8'b00000000;

        map2[16] = 8'b00000000;//3
        map2[17] = 8'b00000000;
        map2[18] = 8'b00000000;
        map2[19] = 8'b00000000;
        map2[20] = 8'b00000000;
        map2[21] = 8'b00000000;
        map2[22] = 8'b00000000;
        map2[23] = 8'b00000000;

        map2[24] = 8'b00000000;//4
        map2[25] = 8'b00000000;
        map2[26] = 8'b00000000;
        map2[27] = 8'b00000000;
        map2[28] = 8'b00000000;
        map2[29] = 8'b00000000;
        map2[30] = 8'b00000000;
        map2[31] = 8'b00000000;

		map2[32] = 8'b00000000;//5
        map2[33] = 8'b00000000;
        map2[34] = 8'b00000000;
        map2[35] = 8'b00000000;
        map2[36] = 8'b00000000;
        map2[37] = 8'b00000000;
        map2[38] = 8'b00000000;
        map2[39] = 8'b00000000;
        
        map2[40] = 8'b00000000;//6
        map2[41] = 8'b00000000;
        map2[42] = 8'b00000000;
        map2[43] = 8'b00000000;
        map2[44] = 8'b00000000;
        map2[45] = 8'b00000000;
        map2[46] = 8'b00000000;
        map2[47] = 8'b00000000;
        
        map2[48] = 8'b00000000;//7
        map2[49] = 8'b00000000;
        map2[50] = 8'b00000000;
        map2[51] = 8'b00000000;
        map2[52] = 8'b00000000;
        map2[53] = 8'b00000000;
        map2[54] = 8'b00000000;
        map2[55] = 8'b00000000;
        
        map2[56] = 8'b00000000;//8
        map2[57] = 8'b00100000;
        map2[58] = 8'b00100000;
        map2[59] = 8'b00100000;
        map2[60] = 8'b00000000;
        map2[61] = 8'b00100000;
        map2[62] = 8'b00000000;
        map2[63] = 8'b00000000;
        
        map2[64] = 8'b00000000;//9
        map2[65] = 8'b00100100;
        map2[66] = 8'b00100100;
        map2[67] = 8'b00100100;
        map2[68] = 8'b00000000;
        map2[69] = 8'b00100100;
        map2[70] = 8'b00000000;
        map2[71] = 8'b00000000;
        
        map2[72] = 8'b00000000;//10
        map2[73] = 8'b00000000;
        map2[74] = 8'b00000000;
        map2[75] = 8'b00000000;
        map2[76] = 8'b00000000;
        map2[77] = 8'b00000000;
        map2[78] = 8'b00000000;
        map2[79] = 8'b00000000;
        
        map2[80] = 8'b01000000;//11
        map2[81] = 8'b00000000;
        map2[82] = 8'b00000000;
        map2[83] = 8'b00000000;
        map2[84] = 8'b00000000;
        map2[85] = 8'b00000000;
        map2[86] = 8'b00000000;
        map2[87] = 8'b00000000;
        
        map2[88] = 8'b00010000;//12
        map2[89] = 8'b00100000;
        map2[90] = 8'b01001000;
        map2[91] = 8'b00000000;
        map2[92] = 8'b00000000;
        map2[93] = 8'b00000000;
        map2[94] = 8'b00000000;
        map2[95] = 8'b00000000;
       
        map2[96] = 8'b00000100;//13
        map2[97] = 8'b00001000;
        map2[98] = 8'b00010000;
        map2[99] = 8'b00100000;
        map2[100] = 8'b01001000;
        map2[101] = 8'b00000000;
        map2[102] = 8'b00000000;
        map2[103] = 8'b00000000;
        
        map2[104] = 8'b00000001;//14
        map2[105] = 8'b00000010;
        map2[106] = 8'b00000100;
        map2[107] = 8'b00001000;
        map2[108] = 8'b10010000;
        map2[109] = 8'b00100000;
        map2[110] = 8'b01000000;
        map2[111] = 8'b10010000;
        
        map2[112] = 8'b00000000;//15
        map2[113] = 8'b00000000;
        map2[114] = 8'b00000001;
        map2[115] = 8'b00000010;
        map2[116] = 8'b00000100;
        map2[117] = 8'b01001000;
        map2[118] = 8'b00010000;
        map2[119] = 8'b00100000;
        
        map2[120] = 8'b00000000;//16
        map2[121] = 8'b00000000;
        map2[122] = 8'b00000000;
        map2[123] = 8'b00000001;
        map2[124] = 8'b00000010;
        map2[125] = 8'b00000100;
        map2[126] = 8'b01001000;
        map2[127] = 8'b00010000;
        
        map2[128] = 8'b00000000;//17
        map2[129] = 8'b00000000;
        map2[130] = 8'b00000000;
        map2[131] = 8'b00000001;
        map2[132] = 8'b00000010;
        map2[133] = 8'b00000100;
        map2[134] = 8'b01001000;
        map2[135] = 8'b00010000;
        
        map2[136] = 8'b00000000;//18
        map2[137] = 8'b00000000;
        map2[138] = 8'b00000000;
        map2[139] = 8'b10000000;
        map2[140] = 8'b10000000;
        map2[141] = 8'b10001001;
        map2[142] = 8'b10000010;
        map2[143] = 8'b00000100;
        
        map2[144] = 8'b00000000;//19
        map2[145] = 8'b00000000;
        map2[146] = 8'b10000000;
        map2[147] = 8'b11000000;
        map2[148] = 8'b01000000;
        map2[149] = 8'b01000000;
        map2[150] = 8'b01010001;
        map2[151] = 8'b10000010;
        
        map2[152] = 8'b00000000;//20
        map2[153] = 8'b00000000;
        map2[154] = 8'b11100000;
        map2[155] = 8'b10110000;
        map2[156] = 8'b00010000;
        map2[157] = 8'b00010000;
        map2[158] = 8'b00010010;
        map2[159] = 8'b10100000;
        
        map2[160] = 8'b00000000;//21
        map2[161] = 8'b00000000;
        map2[162] = 8'b11100000;
        map2[163] = 8'b10110000;
        map2[164] = 8'b00010000;
        map2[165] = 8'b00010000;
        map2[166] = 8'b00010000;
        map2[167] = 8'b10100001;
        
    end
    else
        for(j = 0;j < 168;j = j + 1)
            map2[j] = map2[j];
end

always @(posedge clk or posedge reset_p) begin
    if(reset_p)
    begin
        map3[0] = 8'b00000000;//1
        map3[1] = 8'b00000000;
        map3[2] = 8'b00000000;
        map3[3] = 8'b00000000;
        map3[4] = 8'b10000000;
        map3[5] = 8'b00000000;
        map3[6] = 8'b00000000;
        map3[7] = 8'b00000000;

        map3[8] =  8'b00000000;//2
        map3[9] =  8'b00000000;
        map3[10] = 8'b00000000;
        map3[11] = 8'b10000000;
        map3[12] = 8'b00000000;
        map3[13] = 8'b00000000;
        map3[14] = 8'b00000000;
        map3[15] = 8'b00000000;

        map3[16] = 8'b00000000;//3
        map3[17] = 8'b00000000;
        map3[18] = 8'b00000000;
        map3[19] = 8'b00000000;
        map3[20] = 8'b10000000;
        map3[21] = 8'b00000000;
        map3[22] = 8'b00000000;
        map3[23] = 8'b00000000;

        map3[24] = 8'b00000000;//4
        map3[25] = 8'b00000000;
        map3[26] = 8'b00000000;
        map3[27] = 8'b10000000;
        map3[28] = 8'b00000000;
        map3[29] = 8'b00000000;
        map3[30] = 8'b00000000;
        map3[31] = 8'b00000000;

		map3[32] = 8'b00000000;//5
        map3[33] = 8'b00000000;
        map3[34] = 8'b00000000;
        map3[35] = 8'b00000000;
        map3[36] = 8'b10000000;
        map3[37] = 8'b00000000;
        map3[38] = 8'b00000000;
        map3[39] = 8'b00000000;
        
        map3[40] = 8'b00000000;//6
        map3[41] = 8'b00000000;
        map3[42] = 8'b00000000;
        map3[43] = 8'b00000000;
        map3[44] = 8'b10000000;
        map3[45] = 8'b00000000;
        map3[46] = 8'b00000000;
        map3[47] = 8'b00000000;
        
        map3[48] = 8'b00000000;//7
        map3[49] = 8'b00000000;
        map3[50] = 8'b00000000;
        map3[51] = 8'b00000000;
        map3[52] = 8'b10000000;
        map3[53] = 8'b00000000;
        map3[54] = 8'b00000000;
        map3[55] = 8'b00000000;
        
        map3[56] = 8'b00000000;//8
        map3[57] = 8'b00000000;
        map3[58] = 8'b00000000;
        map3[59] = 8'b00000000;
        map3[60] = 8'b10000000;
        map3[61] = 8'b00000000;
        map3[62] = 8'b00000000;
        map3[63] = 8'b00000000;
        
        map3[64] = 8'b00000000;//9
        map3[65] = 8'b00000000;
        map3[66] = 8'b00000000;
        map3[67] = 8'b00000000;
        map3[68] = 8'b00000000;
        map3[69] = 8'b00000000;
        map3[70] = 8'b00000000;
        map3[71] = 8'b00000000;
        
        map3[72] = 8'b00000000;//10
        map3[73] = 8'b00000000;
        map3[74] = 8'b00000000;
        map3[75] = 8'b00000000;
        map3[76] = 8'b10000000;
        map3[77] = 8'b00000000;
        map3[78] = 8'b00000000;
        map3[79] = 8'b00000000;
        
        map3[80] = 8'b00000000;//11
        map3[81] = 8'b00000000;
        map3[82] = 8'b00000000;
        map3[83] = 8'b00000000;
        map3[84] = 8'b10000000;
        map3[85] = 8'b00000000;
        map3[86] = 8'b00000000;
        map3[87] = 8'b00000000;
        
        map3[88] = 8'b00000000;//12
        map3[89] = 8'b00000000;
        map3[90] = 8'b00000000;
        map3[91] = 8'b00000000;
        map3[92] = 8'b10000000;
        map3[93] = 8'b00000000;
        map3[94] = 8'b00000000;
        map3[95] = 8'b00000000;
       
        map3[96] = 8'b00000000;//13
        map3[97] = 8'b00000000;
        map3[98] = 8'b10000000;
        map3[99] = 8'b00000000;
        map3[100] = 8'b00000000;
        map3[101] = 8'b00000000;
        map3[102] = 8'b10000000;
        map3[103] = 8'b01000000;
        
        map3[104] = 8'b10000000;//14
        map3[105] = 8'b00000000;
        map3[106] = 8'b00000000;
        map3[107] = 8'b00000000;
        map3[108] = 8'b00000000;
        map3[109] = 8'b00000000;
        map3[110] = 8'b10000000;
        map3[111] = 8'b01000000;
        
        map3[112] = 8'b11001000;//15
        map3[113] = 8'b00000000;
        map3[114] = 8'b00000000;
        map3[115] = 8'b00000000;
        map3[116] = 8'b00000000;
        map3[117] = 8'b00000000;
        map3[118] = 8'b10000000;
        map3[119] = 8'b01000000;
        
        map3[120] = 8'b00100000;//16
        map3[121] = 8'b01001000;
        map3[122] = 8'b10000000;
        map3[123] = 8'b00000000;
        map3[124] = 8'b00000000;
        map3[125] = 8'b00000000;
        map3[126] = 8'b10000000;
        map3[127] = 8'b01000000;
        
        map3[128] = 8'b00100000;//17
        map3[129] = 8'b01001000;
        map3[130] = 8'b10000000;
        map3[131] = 8'b00000000;
        map3[132] = 8'b00000000;
        map3[133] = 8'b10000000;
        map3[134] = 8'b10000000;
        map3[135] = 8'b10000000;
        
        map3[136] = 8'b00001000;//18
        map3[137] = 8'b11010010;
        map3[138] = 8'b00000000;
        map3[139] = 8'b00000000;
        map3[140] = 8'b00000000;
        map3[141] = 8'b10000000;
        map3[142] = 8'b10000000;
        map3[143] = 8'b00000000;
        
        map3[144] = 8'b00000100;//19
        map3[145] = 8'b11011000;
        map3[146] = 8'b00100010;
        map3[147] = 8'b00000000;
        map3[148] = 8'b10000000;
        map3[149] = 8'b01000000;
        map3[150] = 8'b10000000;
        map3[151] = 8'b00000000;
        
        map3[152] = 8'b01000000;//20
        map3[153] = 8'b11110111;
        map3[154] = 8'b01001000;
        map3[155] = 8'b11000001;
        map3[156] = 8'b00100000;
        map3[157] = 8'b00100000;
        map3[158] = 8'b01000000;
        map3[159] = 8'b10000000;
        
        map3[160] = 8'b01000000;//21
        map3[161] = 8'b11110111;
        map3[162] = 8'b01001000;
        map3[163] = 8'b11000001;
        map3[164] = 8'b00100000;
        map3[165] = 8'b01000000;
        map3[166] = 8'b10000000;
        map3[167] = 8'b00000000;
        
    end
    else
        for(j = 0;j < 168;j = j + 1)
            map3[j] = map3[j];
end

always @(posedge clk or posedge reset_p) begin
    if(reset_p)
    begin
        map4[0] = 8'b00000000;//1
        map4[1] = 8'b00000000;
        map4[2] = 8'b00000000;
        map4[3] = 8'b00000000;
        map4[4] = 8'b00000000;
        map4[5] = 8'b00000000;
        map4[6] = 8'b00000000;
        map4[7] = 8'b00000000;

        map4[8] = 8'b00000000;//2
        map4[9] = 8'b00000000;
        map4[10] = 8'b00000000;
        map4[11] = 8'b00000000;
        map4[12] = 8'b00000000;
        map4[13] = 8'b00000000;
        map4[14] = 8'b00000000;
        map4[15] = 8'b00000000;

        map4[16] = 8'b00000000;//3
        map4[17] = 8'b00000000;
        map4[18] = 8'b00000000;
        map4[19] = 8'b00000000;
        map4[20] = 8'b00000000;
        map4[21] = 8'b00000000;
        map4[22] = 8'b00000000;
        map4[23] = 8'b00000000;

        map4[24] = 8'b00000000;//4
        map4[25] = 8'b00000000;
        map4[26] = 8'b00000000;
        map4[27] = 8'b00000000;
        map4[28] = 8'b00000000;
        map4[29] = 8'b00000000;
        map4[30] = 8'b00000000;
        map4[31] = 8'b00000000;

		map4[32] = 8'b00000000;//5
        map4[33] = 8'b00000000;
        map4[34] = 8'b00000000;
        map4[35] = 8'b00000000;
        map4[36] = 8'b00000000;
        map4[37] = 8'b00000000;
        map4[38] = 8'b00000000;
        map4[39] = 8'b00000000;
        
        map4[40] = 8'b00000000;//6
        map4[41] = 8'b00000000;
        map4[42] = 8'b00000000;
        map4[43] = 8'b00000000;
        map4[44] = 8'b00000000;
        map4[45] = 8'b00000000;
        map4[46] = 8'b00000000;
        map4[47] = 8'b00000000;
        
        map4[48] = 8'b00000000;//7
        map4[49] = 8'b00000000;
        map4[50] = 8'b00000000;
        map4[51] = 8'b00000000;
        map4[52] = 8'b00000000;
        map4[53] = 8'b00000000;
        map4[54] = 8'b00000000;
        map4[55] = 8'b00000000;
        
        map4[56] = 8'b00000000;//8
        map4[57] = 8'b00000000;
        map4[58] = 8'b00000000;
        map4[59] = 8'b00000000;
        map4[60] = 8'b00000000;
        map4[61] = 8'b00000000;
        map4[62] = 8'b00000000;
        map4[63] = 8'b00000000;
        
        map4[64] = 8'b00000000;//9
        map4[65] = 8'b00000000;
        map4[66] = 8'b00000000;
        map4[67] = 8'b00000000;
        map4[68] = 8'b00000000;
        map4[69] = 8'b00000000;
        map4[70] = 8'b00000000;
        map4[71] = 8'b00000000;
        
        map4[72] = 8'b00000000;//10
        map4[73] = 8'b00000000;
        map4[74] = 8'b00000000;
        map4[75] = 8'b00000000;
        map4[76] = 8'b00000000;
        map4[77] = 8'b00000000;
        map4[78] = 8'b00000000;
        map4[79] = 8'b00000000;
        
        map4[80] = 8'b00000000;//11
        map4[81] = 8'b00000000;
        map4[82] = 8'b00000000;
        map4[83] = 8'b00000000;
        map4[84] = 8'b00000000;
        map4[85] = 8'b00000000;
        map4[86] = 8'b00000000;
        map4[87] = 8'b00000000;
        
        map4[88] = 8'b00000000;//12
        map4[89] = 8'b00000000;
        map4[90] = 8'b00000000;
        map4[91] = 8'b00000000;
        map4[92] = 8'b00000000;
        map4[93] = 8'b00000000;
        map4[94] = 8'b00000000;
        map4[95] = 8'b00000000;
       
        map4[96] =  8'b00000000;//13
        map4[97] =  8'b00000000;
        map4[98] =  8'b00000000;
        map4[99] =  8'b00000001;
        map4[100] = 8'b00000001;
        map4[101] = 8'b00000010;
        map4[102] = 8'b00000010;
        map4[103] = 8'b00000010;
        
        map4[104] = 8'b00000000;//14
        map4[105] = 8'b00000000;
        map4[106] = 8'b00000001;
        map4[107] = 8'b00000010;
        map4[108] = 8'b00000010;
        map4[109] = 8'b00000100;
        map4[110] = 8'b00000100;
        map4[111] = 8'b00000101;
        
        map4[112] = 8'b00000000;//15
        map4[113] = 8'b00000001;
        map4[114] = 8'b10000010;
        map4[115] = 8'b00000100;
        map4[116] = 8'b00000100;
        map4[117] = 8'b00001000;
        map4[118] = 8'b00001001;
        map4[119] = 8'b00001010;
        
        map4[120] = 8'b00000000;//16
        map4[121] = 8'b00000000;
        map4[122] = 8'b00000010;
        map4[123] = 8'b10000101;
        map4[124] = 8'b00001000;
        map4[125] = 8'b00001000;
        map4[126] = 8'b00010000;
        map4[127] = 8'b00010010;
        
        map4[128] = 8'b00000000;//17
        map4[129] = 8'b00000000;
        map4[130] = 8'b00000010;
        map4[131] = 8'b00000101;
        map4[132] = 8'b00001000;
        map4[133] = 8'b00001000;
        map4[134] = 8'b00010000;
        map4[135] = 8'b00010010;
        
        map4[136] = 8'b00000000;//18
        map4[137] = 8'b00000000;
        map4[138] = 8'b00000010;
        map4[139] = 8'b01000101;
        map4[140] = 8'b10001000;
        map4[141] = 8'b00001000;
        map4[142] = 8'b00010000;
        map4[143] = 8'b00010010;
        
        map4[144] = 8'b00000000;//19
        map4[145] = 8'b00000000;
        map4[146] = 8'b00000010;
        map4[147] = 8'b00000101;
        map4[148] = 8'b01001000;
        map4[149] = 8'b10001000;
        map4[150] = 8'b00010000;
        map4[151] = 8'b00010010;
        
        map4[152] = 8'b00000000;//20
        map4[153] = 8'b00000000;
        map4[154] = 8'b00000010;
        map4[155] = 8'b00000101;
        map4[156] = 8'b00001000;
        map4[157] = 8'b00001000;
        map4[158] = 8'b00110000;
        map4[159] = 8'b01010010;
        
        map4[160] = 8'b00000000;//21
        map4[161] = 8'b00000000;
        map4[162] = 8'b00000010;
        map4[163] = 8'b00000101;
        map4[164] = 8'b00001000;
        map4[165] = 8'b00001000;
        map4[166] = 8'b00010000;
        map4[167] = 8'b00110010;
        
    end
    else
        for(j = 0;j < 168;j = j + 1)
            map4[j] = map4[j];
end
/*
always @(posedge clk or posedge reset_p) begin
    if(reset_p)
    begin
        map[0] = 8'b00000000;//1
        map[1] = 8'b00000000;
        map[2] = 8'b00000000;
        map[3] = 8'b00000000;
        map[4] = 8'b00000000;
        map[5] = 8'b00000000;
        map[6] = 8'b00000000;
        map[7] = 8'b00000000;

        map[8] = 8'b00000000;//2
        map[9] = 8'b00000000;
        map[10] = 8'b00000000;
        map[11] = 8'b00000000;
        map[12] = 8'b00000000;
        map[13] = 8'b00000000;
        map[14] = 8'b00000000;
        map[15] = 8'b00000000;

        map[16] = 8'b00000000;//3
        map[17] = 8'b00000000;
        map[18] = 8'b00000000;
        map[19] = 8'b00000000;
        map[20] = 8'b00000000;
        map[21] = 8'b00000000;
        map[22] = 8'b00000000;
        map[23] = 8'b00000000;

        map[24] = 8'b00000000;//4
        map[25] = 8'b00000000;
        map[26] = 8'b00000000;
        map[27] = 8'b00000000;
        map[28] = 8'b00000000;
        map[29] = 8'b00000000;
        map[30] = 8'b00000000;
        map[31] = 8'b00000000;

		map[32] = 8'b00000000;//5
        map[33] = 8'b00000000;
        map[34] = 8'b00000000;
        map[35] = 8'b00000000;
        map[36] = 8'b00000000;
        map[37] = 8'b00000000;
        map[38] = 8'b00000000;
        map[39] = 8'b00000000;
        
        map[40] = 8'b00000000;//6
        map[41] = 8'b00000000;
        map[42] = 8'b00000000;
        map[43] = 8'b00000000;
        map[44] = 8'b00000000;
        map[45] = 8'b00000000;
        map[46] = 8'b00000000;
        map[47] = 8'b00000000;
        
        map[48] = 8'b00000000;//7
        map[49] = 8'b00000000;
        map[50] = 8'b00000000;
        map[51] = 8'b00000000;
        map[52] = 8'b00000000;
        map[53] = 8'b00000000;
        map[54] = 8'b00000000;
        map[55] = 8'b00000000;
        
        map[56] = 8'b00000000;//8
        map[57] = 8'b00000000;
        map[58] = 8'b00000000;
        map[59] = 8'b00000000;
        map[60] = 8'b00000000;
        map[61] = 8'b00000000;
        map[62] = 8'b00000000;
        map[63] = 8'b00000000;
        
        map[64] = 8'b00000000;//9
        map[65] = 8'b00000000;
        map[66] = 8'b00000000;
        map[67] = 8'b00000000;
        map[68] = 8'b00000000;
        map[69] = 8'b00000000;
        map[70] = 8'b00000000;
        map[71] = 8'b00000000;
        
        map[72] = 8'b00000000;//10
        map[73] = 8'b00000000;
        map[74] = 8'b00000000;
        map[75] = 8'b00000000;
        map[76] = 8'b00000000;
        map[77] = 8'b00000000;
        map[78] = 8'b00000000;
        map[79] = 8'b00000000;
        
        map[80] = 8'b00000000;//11
        map[81] = 8'b00000000;
        map[82] = 8'b00000000;
        map[83] = 8'b00000000;
        map[84] = 8'b00000000;
        map[85] = 8'b00000000;
        map[86] = 8'b00000000;
        map[87] = 8'b00000000;
        
        map[88] = 8'b00000000;//12
        map[89] = 8'b00000000;
        map[90] = 8'b00000000;
        map[91] = 8'b00000000;
        map[92] = 8'b00000000;
        map[93] = 8'b00000000;
        map[94] = 8'b00000000;
        map[95] = 8'b00000000;
       
        map[96] = 8'b00000000;//13
        map[97] = 8'b00000000;
        map[98] = 8'b00000000;
        map[99] = 8'b00000000;
        map[100] = 8'b00000000;
        map[101] = 8'b00000000;
        map[102] = 8'b00000000;
        map[103] = 8'b00000000;
        
        map[104] = 8'b00000000;//14
        map[105] = 8'b00000000;
        map[106] = 8'b00000000;
        map[107] = 8'b00000000;
        map[108] = 8'b00000000;
        map[109] = 8'b00000000;
        map[110] = 8'b00000000;
        map[111] = 8'b00000000;
        
        map[112] = 8'b00000000;//15
        map[113] = 8'b00000000;
        map[114] = 8'b00000000;
        map[115] = 8'b00000000;
        map[116] = 8'b00000000;
        map[117] = 8'b00000000;
        map[118] = 8'b00000000;
        map[119] = 8'b00000000;
        
        map[120] = 8'b00000000;//16
        map[121] = 8'b00000000;
        map[122] = 8'b00000000;
        map[123] = 8'b00000000;
        map[124] = 8'b00000000;
        map[125] = 8'b00000000;
        map[126] = 8'b00000000;
        map[127] = 8'b00000000;
        
        map[128] = 8'b00000000;//17
        map[129] = 8'b00000000;
        map[130] = 8'b00000000;
        map[131] = 8'b00000000;
        map[132] = 8'b00000000;
        map[133] = 8'b00000000;
        map[134] = 8'b00000000;
        map[135] = 8'b00000000;
        
        map[136] = 8'b00000000;//18
        map[137] = 8'b00000000;
        map[138] = 8'b00000000;
        map[139] = 8'b00000000;
        map[140] = 8'b00000000;
        map[141] = 8'b00000000;
        map[142] = 8'b00000000;
        map[143] = 8'b00000000;
        
        map[144] = 8'b00000000;//19
        map[145] = 8'b00000000;
        map[146] = 8'b00000000;
        map[147] = 8'b00000000;
        map[148] = 8'b00000000;
        map[149] = 8'b00000000;
        map[150] = 8'b00000000;
        map[151] = 8'b00000000;
        
        map[152] = 8'b00000000;//20
        map[153] = 8'b00000000;
        map[154] = 8'b00000000;
        map[155] = 8'b00000000;
        map[156] = 8'b00000000;
        map[157] = 8'b00000000;
        map[158] = 8'b00000000;
        map[159] = 8'b00000000;
        
        map[160] = 8'b00000000;//21
        map[161] = 8'b00000000;
        map[162] = 8'b00000000;
        map[163] = 8'b00000000;
        map[164] = 8'b00000000;
        map[165] = 8'b00000000;
        map[166] = 8'b00000000;
        map[167] = 8'b00000000;
        
    end
    else
        for(j = 0;j < 168;j = j + 1)
            map[j] = map[j];
end
always @(posedge clk or posedge reset_p) begin
    if(reset_p)
    begin
        map[0] = 8'b00000000;//1
        map[1] = 8'b00000000;
        map[2] = 8'b00000000;
        map[3] = 8'b00000000;
        map[4] = 8'b00000000;
        map[5] = 8'b00000000;
        map[6] = 8'b00000000;
        map[7] = 8'b00000000;

        map[8] = 8'b00000000;//2
        map[9] = 8'b00000000;
        map[10] = 8'b00000000;
        map[11] = 8'b00000000;
        map[12] = 8'b00000000;
        map[13] = 8'b00000000;
        map[14] = 8'b00000000;
        map[15] = 8'b00000000;

        map[16] = 8'b00000000;//3
        map[17] = 8'b00000000;
        map[18] = 8'b00000000;
        map[19] = 8'b00000000;
        map[20] = 8'b00000000;
        map[21] = 8'b00000000;
        map[22] = 8'b00000000;
        map[23] = 8'b00000000;

        map[24] = 8'b00000000;//4
        map[25] = 8'b00000000;
        map[26] = 8'b00000000;
        map[27] = 8'b00000000;
        map[28] = 8'b00000000;
        map[29] = 8'b00000000;
        map[30] = 8'b00000000;
        map[31] = 8'b00000000;

		map[32] = 8'b00000000;//5
        map[33] = 8'b00000000;
        map[34] = 8'b00000000;
        map[35] = 8'b00000000;
        map[36] = 8'b00000000;
        map[37] = 8'b00000000;
        map[38] = 8'b00000000;
        map[39] = 8'b00000000;
        
        map[40] = 8'b00000000;//6
        map[41] = 8'b00000000;
        map[42] = 8'b00000000;
        map[43] = 8'b00000000;
        map[44] = 8'b00000000;
        map[45] = 8'b00000000;
        map[46] = 8'b00000000;
        map[47] = 8'b00000000;
        
        map[48] = 8'b00000000;//7
        map[49] = 8'b00000000;
        map[50] = 8'b00000000;
        map[51] = 8'b00000000;
        map[52] = 8'b00000000;
        map[53] = 8'b00000000;
        map[54] = 8'b00000000;
        map[55] = 8'b00000000;
        
        map[56] = 8'b00000000;//8
        map[57] = 8'b00000000;
        map[58] = 8'b00000000;
        map[59] = 8'b00000000;
        map[60] = 8'b00000000;
        map[61] = 8'b00000000;
        map[62] = 8'b00000000;
        map[63] = 8'b00000000;
        
        map[64] = 8'b00000000;//9
        map[65] = 8'b00000000;
        map[66] = 8'b00000000;
        map[67] = 8'b00000000;
        map[68] = 8'b00000000;
        map[69] = 8'b00000000;
        map[70] = 8'b00000000;
        map[71] = 8'b00000000;
        
        map[72] = 8'b00000000;//10
        map[73] = 8'b00000000;
        map[74] = 8'b00000000;
        map[75] = 8'b00000000;
        map[76] = 8'b00000000;
        map[77] = 8'b00000000;
        map[78] = 8'b00000000;
        map[79] = 8'b00000000;
        
        map[80] = 8'b00000000;//11
        map[81] = 8'b00000000;
        map[82] = 8'b00000000;
        map[83] = 8'b00000000;
        map[84] = 8'b00000000;
        map[85] = 8'b00000000;
        map[86] = 8'b00000000;
        map[87] = 8'b00000000;
        
        map[88] = 8'b00000000;//12
        map[89] = 8'b00000000;
        map[90] = 8'b00000000;
        map[91] = 8'b00000000;
        map[92] = 8'b00000000;
        map[93] = 8'b00000000;
        map[94] = 8'b00000000;
        map[95] = 8'b00000000;
       
        map[96] = 8'b00000000;//13
        map[97] = 8'b00000000;
        map[98] = 8'b00000000;
        map[99] = 8'b00000000;
        map[100] = 8'b00000000;
        map[101] = 8'b00000000;
        map[102] = 8'b00000000;
        map[103] = 8'b00000000;
        
        map[104] = 8'b00000000;//14
        map[105] = 8'b00000000;
        map[106] = 8'b00000000;
        map[107] = 8'b00000000;
        map[108] = 8'b00000000;
        map[109] = 8'b00000000;
        map[110] = 8'b00000000;
        map[111] = 8'b00000000;
        
        map[112] = 8'b00000000;//15
        map[113] = 8'b00000000;
        map[114] = 8'b00000000;
        map[115] = 8'b00000000;
        map[116] = 8'b00000000;
        map[117] = 8'b00000000;
        map[118] = 8'b00000000;
        map[119] = 8'b00000000;
        
        map[120] = 8'b00000000;//16
        map[121] = 8'b00000000;
        map[122] = 8'b00000000;
        map[123] = 8'b00000000;
        map[124] = 8'b00000000;
        map[125] = 8'b00000000;
        map[126] = 8'b00000000;
        map[127] = 8'b00000000;
        
        map[128] = 8'b00000000;//17
        map[129] = 8'b00000000;
        map[130] = 8'b00000000;
        map[131] = 8'b00000000;
        map[132] = 8'b00000000;
        map[133] = 8'b00000000;
        map[134] = 8'b00000000;
        map[135] = 8'b00000000;
        
        map[136] = 8'b00000000;//18
        map[137] = 8'b00000000;
        map[138] = 8'b00000000;
        map[139] = 8'b00000000;
        map[140] = 8'b00000000;
        map[141] = 8'b00000000;
        map[142] = 8'b00000000;
        map[143] = 8'b00000000;
        
        map[144] = 8'b00000000;//19
        map[145] = 8'b00000000;
        map[146] = 8'b00000000;
        map[147] = 8'b00000000;
        map[148] = 8'b00000000;
        map[149] = 8'b00000000;
        map[150] = 8'b00000000;
        map[151] = 8'b00000000;
        
        map[152] = 8'b00000000;//20
        map[153] = 8'b00000000;
        map[154] = 8'b00000000;
        map[155] = 8'b00000000;
        map[156] = 8'b00000000;
        map[157] = 8'b00000000;
        map[158] = 8'b00000000;
        map[159] = 8'b00000000;
        
        map[160] = 8'b00000000;//21
        map[161] = 8'b00000000;
        map[162] = 8'b00000000;
        map[163] = 8'b00000000;
        map[164] = 8'b00000000;
        map[165] = 8'b00000000;
        map[166] = 8'b00000000;
        map[167] = 8'b00000000;
        
    end
    else
        for(j = 0;j < 168;j = j + 1)
            map[j] = map[j];
end
always @(posedge clk or posedge reset_p) begin
    if(reset_p)
    begin
        map[0] = 8'b00000000;//1
        map[1] = 8'b00000000;
        map[2] = 8'b00000000;
        map[3] = 8'b00000000;
        map[4] = 8'b00000000;
        map[5] = 8'b00000000;
        map[6] = 8'b00000000;
        map[7] = 8'b00000000;

        map[8] = 8'b00000000;//2
        map[9] = 8'b00000000;
        map[10] = 8'b00000000;
        map[11] = 8'b00000000;
        map[12] = 8'b00000000;
        map[13] = 8'b00000000;
        map[14] = 8'b00000000;
        map[15] = 8'b00000000;

        map[16] = 8'b00000000;//3
        map[17] = 8'b00000000;
        map[18] = 8'b00000000;
        map[19] = 8'b00000000;
        map[20] = 8'b00000000;
        map[21] = 8'b00000000;
        map[22] = 8'b00000000;
        map[23] = 8'b00000000;

        map[24] = 8'b00000000;//4
        map[25] = 8'b00000000;
        map[26] = 8'b00000000;
        map[27] = 8'b00000000;
        map[28] = 8'b00000000;
        map[29] = 8'b00000000;
        map[30] = 8'b00000000;
        map[31] = 8'b00000000;

		map[32] = 8'b00000000;//5
        map[33] = 8'b00000000;
        map[34] = 8'b00000000;
        map[35] = 8'b00000000;
        map[36] = 8'b00000000;
        map[37] = 8'b00000000;
        map[38] = 8'b00000000;
        map[39] = 8'b00000000;
        
        map[40] = 8'b00000000;//6
        map[41] = 8'b00000000;
        map[42] = 8'b00000000;
        map[43] = 8'b00000000;
        map[44] = 8'b00000000;
        map[45] = 8'b00000000;
        map[46] = 8'b00000000;
        map[47] = 8'b00000000;
        
        map[48] = 8'b00000000;//7
        map[49] = 8'b00000000;
        map[50] = 8'b00000000;
        map[51] = 8'b00000000;
        map[52] = 8'b00000000;
        map[53] = 8'b00000000;
        map[54] = 8'b00000000;
        map[55] = 8'b00000000;
        
        map[56] = 8'b00000000;//8
        map[57] = 8'b00000000;
        map[58] = 8'b00000000;
        map[59] = 8'b00000000;
        map[60] = 8'b00000000;
        map[61] = 8'b00000000;
        map[62] = 8'b00000000;
        map[63] = 8'b00000000;
        
        map[64] = 8'b00000000;//9
        map[65] = 8'b00000000;
        map[66] = 8'b00000000;
        map[67] = 8'b00000000;
        map[68] = 8'b00000000;
        map[69] = 8'b00000000;
        map[70] = 8'b00000000;
        map[71] = 8'b00000000;
        
        map[72] = 8'b00000000;//10
        map[73] = 8'b00000000;
        map[74] = 8'b00000000;
        map[75] = 8'b00000000;
        map[76] = 8'b00000000;
        map[77] = 8'b00000000;
        map[78] = 8'b00000000;
        map[79] = 8'b00000000;
        
        map[80] = 8'b00000000;//11
        map[81] = 8'b00000000;
        map[82] = 8'b00000000;
        map[83] = 8'b00000000;
        map[84] = 8'b00000000;
        map[85] = 8'b00000000;
        map[86] = 8'b00000000;
        map[87] = 8'b00000000;
        
        map[88] = 8'b00000000;//12
        map[89] = 8'b00000000;
        map[90] = 8'b00000000;
        map[91] = 8'b00000000;
        map[92] = 8'b00000000;
        map[93] = 8'b00000000;
        map[94] = 8'b00000000;
        map[95] = 8'b00000000;
       
        map[96] = 8'b00000000;//13
        map[97] = 8'b00000000;
        map[98] = 8'b00000000;
        map[99] = 8'b00000000;
        map[100] = 8'b00000000;
        map[101] = 8'b00000000;
        map[102] = 8'b00000000;
        map[103] = 8'b00000000;
        
        map[104] = 8'b00000000;//14
        map[105] = 8'b00000000;
        map[106] = 8'b00000000;
        map[107] = 8'b00000000;
        map[108] = 8'b00000000;
        map[109] = 8'b00000000;
        map[110] = 8'b00000000;
        map[111] = 8'b00000000;
        
        map[112] = 8'b00000000;//15
        map[113] = 8'b00000000;
        map[114] = 8'b00000000;
        map[115] = 8'b00000000;
        map[116] = 8'b00000000;
        map[117] = 8'b00000000;
        map[118] = 8'b00000000;
        map[119] = 8'b00000000;
        
        map[120] = 8'b00000000;//16
        map[121] = 8'b00000000;
        map[122] = 8'b00000000;
        map[123] = 8'b00000000;
        map[124] = 8'b00000000;
        map[125] = 8'b00000000;
        map[126] = 8'b00000000;
        map[127] = 8'b00000000;
        
        map[128] = 8'b00000000;//17
        map[129] = 8'b00000000;
        map[130] = 8'b00000000;
        map[131] = 8'b00000000;
        map[132] = 8'b00000000;
        map[133] = 8'b00000000;
        map[134] = 8'b00000000;
        map[135] = 8'b00000000;
        
        map[136] = 8'b00000000;//18
        map[137] = 8'b00000000;
        map[138] = 8'b00000000;
        map[139] = 8'b00000000;
        map[140] = 8'b00000000;
        map[141] = 8'b00000000;
        map[142] = 8'b00000000;
        map[143] = 8'b00000000;
        
        map[144] = 8'b00000000;//19
        map[145] = 8'b00000000;
        map[146] = 8'b00000000;
        map[147] = 8'b00000000;
        map[148] = 8'b00000000;
        map[149] = 8'b00000000;
        map[150] = 8'b00000000;
        map[151] = 8'b00000000;
        
        map[152] = 8'b00000000;//20
        map[153] = 8'b00000000;
        map[154] = 8'b00000000;
        map[155] = 8'b00000000;
        map[156] = 8'b00000000;
        map[157] = 8'b00000000;
        map[158] = 8'b00000000;
        map[159] = 8'b00000000;
        
        map[160] = 8'b00000000;//21
        map[161] = 8'b00000000;
        map[162] = 8'b00000000;
        map[163] = 8'b00000000;
        map[164] = 8'b00000000;
        map[165] = 8'b00000000;
        map[166] = 8'b00000000;
        map[167] = 8'b00000000;
        
    end
    else
        for(j = 0;j < 168;j = j + 1)
            map[j] = map[j];
end*/

endmodule